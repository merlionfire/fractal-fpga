parameter     REG_MOUSE_CTRL_STATUS_ADDR   = 4'h0 ;
parameter     REG_CURSOR_COLOR_ADDR        = 4'h4 ;
parameter     REG_CURSOR_X_LOW_ADDR        = 4'h5 ;
parameter     REG_CURSOR_X_HIGH_ADDR       = 4'h6 ;
parameter     REG_CURSOR_Y_LOW_ADDR        = 4'h7 ;
parameter     REG_CURSOR_Y_HIGH_ADDR       = 4'h8 ;
parameter     REG_SEL_X_LEFT_LOW_ADDR      = 4'h9 ; 
parameter     REG_SEL_X_LEFT_HIGH_ADDR     = 4'hA ;
parameter     REG_SEL_Y_BOT_LOW_ADDR       = 4'hB ;
parameter     REG_SEL_Y_BOT_HIGH_ADDR      = 4'hC ; 
parameter     REG_SEL_HALF_LENGTH_LOW_ADDR      = 4'hE ;
parameter     REG_SEL_HALF_LENGTH_HIGH_ADDR     = 4'hF ;

