
 parameter  REG_ALU_CTRL_STATUS_ADDR      =  4'h0;
 parameter  REG_ALU_A_0_ADDR              =  4'h1;
 parameter  REG_ALU_A_1_ADDR              =  4'h2;
 parameter  REG_ALU_A_2_ADDR              =  4'h3;
 parameter  REG_ALU_A_3_ADDR              =  4'h4;
 parameter  REG_ALU_B_0_ADDR              =  4'h5;
 parameter  REG_ALU_B_1_ADDR              =  4'h6;
 parameter  REG_ALU_B_2_ADDR              =  4'h7;
 parameter  REG_ALU_B_3_ADDR              =  4'h8;
 parameter  REG_ALU_Q_0_ADDR              =  4'h1;
 parameter  REG_ALU_Q_1_ADDR              =  4'h2;
 parameter  REG_ALU_Q_2_ADDR              =  4'h3;
 parameter  REG_ALU_Q_3_ADDR              =  4'h4;
 parameter  REG_ALU_R_0_ADDR              =  4'h5;
 parameter  REG_ALU_R_1_ADDR              =  4'h6;
 parameter  REG_ALU_R_2_ADDR              =  4'h7;
 parameter  REG_ALU_R_3_ADDR              =  4'h8;
