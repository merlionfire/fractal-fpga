

module char_buffer_wrapper (
   input  wire        clk,
   input  wire [10:0] cb_rd_addr,
   output wire [7:0]  cb_rd_data,
   input  wire [10:0] cb_wr_addr,
   input  wire        cb_wr_en,
   input  wire [7:0]  cb_wr_data
); 


//   number of chars 
// = (pixel_x / font_width_pixel ) * ( pixel_y / font_height_pixel ) 
// = ( 1024 / 8 ) X ( 768 / 16 ) 
// = 128 X 48 
// = 6 * 1024 = 6K bytes  

   RAMB16_S9_S9 #(
    .INIT_A  ( 9'h020 ),     
    .INIT_B  ( 9'h020 ),     
    .INIT_00 ( 256'h30_30_40_5A_59_58_57_56_55_54_53_52_51_50_4F_4E_4D_4C_4B_4A_49_48_47_46_45_44_43_42_41_40_30_30 ),
    .INIT_01 ( 256'h31_30_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_31_30 ),
    .INIT_02 ( 256'h32_30_20_20_20_20_4C_41_54_43_41_52_46_20_54_45_53_20_54_4F_52_42_4C_45_44_4E_41_4D_20_20_32_30 ),
    .INIT_03 ( 256'h33_30_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_33_30 ),
    .INIT_04 ( 256'h34_30_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_3A_52_45_54_45_4D_41_52_41_50_20_34_30 ),
    .INIT_05 ( 256'h35_30_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_3A_78_20_20_20_74_66_65_6C_20_2D_20_35_30 ),
    .INIT_06 ( 256'h36_30_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_3A_79_20_6D_6F_74_74_6F_62_20_2D_20_36_30 ),
    .INIT_07 ( 256'h37_30_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_3A_20_20_20_61_74_6C_65_64_20_2D_20_37_30 ),
    .INIT_08 ( 256'h38_30_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_3A_72_65_74_69_20_78_61_6D_20_2D_20_38_30 ),
    .INIT_09 ( 256'h39_30_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_39_30 ),
    .INIT_0A ( 256'h30_31_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_30_31 ),
    .INIT_0B ( 256'h31_31_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_3A_50_4C_45_48_20_31_31 ),
    .INIT_0C ( 256'h32_31_20_20_74_65_73_20_6F_74_20_65_73_75_6F_6D_20_73_73_65_72_70_20_74_66_65_4C_20_2D_20_32_31 ),
    .INIT_0D ( 256'h33_31_20_20_20_20_2E_6E_6F_69_67_65_72_20_77_65_6E_20_66_6F_20_72_65_74_6E_65_63_20_20_20_33_31 ),
    .INIT_0E ( 256'h34_31_20_20_20_6F_74_20_65_73_75_6F_6D_20_65_76_6F_6D_20_64_6E_61_20_64_6C_6F_48_20_20_20_34_31 ),
    .INIT_0F ( 256'h35_31_20_20_20_20_20_20_20_20_20_20_20_2E_6E_6F_69_67_65_72_20_74_63_65_6C_65_73_20_20_20_35_31 ),
    .INIT_10 ( 256'h36_31_20_20_20_20_77_61_72_64_20_6F_74_20_65_73_75_6F_6D_20_65_73_61_65_6C_65_52_20_20_20_36_31 ),
    .INIT_11 ( 256'h37_31_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_2E_65_67_61_6D_69_20_77_65_6E_20_20_20_37_31 ),
    .INIT_12 ( 256'h38_31_20_20_20_20_20_6F_74_20_65_73_75_6F_6D_20_6B_63_69_6C_63_20_74_68_67_69_52_20_2D_20_38_31 ),
    .INIT_13 ( 256'h39_31_20_20_20_2E_65_67_61_6D_69_20_6C_61_69_74_69_6E_69_20_65_72_6F_74_73_65_72_20_20_20_39_31 ),
    .INIT_14 ( 256'h30_32_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_30_32 ),
    .INIT_15 ( 256'h31_32_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_31_32 ),
    .INIT_16 ( 256'h32_32_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_32_32 ),
    .INIT_17 ( 256'h33_32_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_33_32 ),
    .INIT_18 ( 256'h34_32_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_34_32 ),
    .INIT_19 ( 256'h35_32_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_35_32 ),
    .INIT_1A ( 256'h36_32_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_36_32 ),
    .INIT_1B ( 256'h37_32_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_37_32 ),
    .INIT_1C ( 256'h38_32_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_38_32 ),
    .INIT_1D ( 256'h39_32_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_39_32 ),
    .INIT_1E ( 256'h30_33_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_30_33 ),
    .INIT_1F ( 256'h31_33_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_31_33 ),
    .INIT_20 ( 256'h32_33_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_32_33 ),
    .INIT_21 ( 256'h33_33_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_33_33 ),
    .INIT_22 ( 256'h34_33_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_34_33 ),
    .INIT_23 ( 256'h35_33_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_35_33 ),
    .INIT_24 ( 256'h36_33_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_36_33 ),
    .INIT_25 ( 256'h37_33_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_37_33 ),
    .INIT_26 ( 256'h38_33_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_38_33 ),
    .INIT_27 ( 256'h39_33_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_39_33 ),
    .INIT_28 ( 256'h30_34_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_30_34 ),
    .INIT_29 ( 256'h31_34_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_31_34 ),
    .INIT_2A ( 256'h32_34_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_32_34 ),
    .INIT_2B ( 256'h33_34_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_33_34 ),
    .INIT_2C ( 256'h34_34_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_34_34 ),
    .INIT_2D ( 256'h35_34_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_35_34 ),
    .INIT_2E ( 256'h36_34_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_36_34 ),
    .INIT_2F ( 256'h37_34_40_5A_59_58_57_56_55_54_53_52_51_50_4F_4E_4D_4C_4B_4A_49_48_47_46_45_44_43_42_41_40_37_34 ),
    .INIT_30 ( 256'h38_34_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_38_34 ),
    .INIT_31 ( 256'h39_34_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_39_34 ),
    .INIT_32 ( 256'h30_35_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_30_35 ),
    .INIT_33 ( 256'h31_35_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_31_35 ),
    .INIT_34 ( 256'h32_35_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_32_35 ),
    .INIT_35 ( 256'h33_35_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_33_35 ),
    .INIT_36 ( 256'h34_35_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_34_35 ),
    .INIT_37 ( 256'h35_35_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_35_35 ),
    .INIT_38 ( 256'h36_35_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_36_35 ),
    .INIT_39 ( 256'h37_35_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_37_35 ),
    .INIT_3A ( 256'h38_35_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_38_35 ),
    .INIT_3B ( 256'h39_35_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_39_35 ),
    .INIT_3C ( 256'h30_36_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_30_36 ),
    .INIT_3D ( 256'h31_36_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_31_36 ),
    .INIT_3E ( 256'h32_36_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_32_36 ),
    .INIT_3F ( 256'h33_36_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_20_33_36 ),
    .SIM_COLLISION_CHECK("NONE")
   ) char_buffer_inst (
    .CLKA   ( clk        ),
    .ADDRA  ( cb_rd_addr ),
    .ENA    ( 1'b1       ),
    .DIA    ( 8'h00      ),
    .DIPA   ( 1'b0       ),
    .WEA    ( 1'b0       ),
    .DOA    ( cb_rd_data ),
    .DOPA   (            ),
    .SSRA   ( 1'b0       ),
    .CLKB   ( clk        ),
    .ADDRB  ( cb_wr_addr ),
    .ENB    ( 1'b1       ),
    .DIB    ( cb_wr_data ),
    .DIPB   ( 1'b0       ),
    .WEB    ( cb_wr_en   ),
    .DOB    (            ),
    .DOPB   (            ),
    .SSRB   ( 1'b0       )
   );

endmodule 
