package env_pkg;
   import uvm_pkg::*;
   import stimulus_pkg::*;

   `include "driver.sv"
   `include "write_monitor.sv"
   `include "master_agent.sv"
   `include "reset_driver.sv"
   `include "reset_agent.sv"
   `include "reset_monitor.sv"
   `include "read_monitor.sv"
   `include "output_agent.sv"
   `include "scoreboard.sv"
   `include "fractal_env.sv"

endpackage 
