package  stimulus_pkg;
   import uvm_pkg::*;
   `include "packet.sv" 
   `include "packet_sequence.sv"
   `include "ports_reset_sequence.sv"
   `include "reset_tr.sv"
   `include "reset_sequence.sv"
   `include "virtual_reset_sequence.sv"
   `include "transformer.sv"
endpackage 
