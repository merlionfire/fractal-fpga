`include "test_base.sv"
