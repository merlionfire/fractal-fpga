`define MAX_SEL_NUM  17
