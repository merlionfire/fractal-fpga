
parameter   REG_CW_CS_ADDR                   =  4'h0; 
parameter   REG_CW_X_ORIG_ADDR               =  4'h1;
parameter   REG_CW_Y_ORIG_ADDR               =  4'h2;
parameter   REG_CW_X_SIZE_ADDR               =  4'h3;
parameter   REG_CW_Y_SIZE_ADDR               =  4'h4;
parameter   REG_CB_ADDR_ORIG_LOW_ADDR        =  4'h5; 
parameter   REG_CB_ADDR_ORIG_HIGH_ADDR       =  4'h6;
parameter   REG_CHAR_RGL_ADDR                =  4'h7;
parameter   REG_GRAPH_BG_RGL_ADDR            =  4'h8;
parameter   REG_CW_ROW_ADDR                  =  4'h9;
parameter   REG_CW_COL_ADDR                  =  4'ha;
parameter   REG_CB_WR_DATA                   =  4'hb;
