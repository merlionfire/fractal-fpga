parameter REG_UART_STATUS_ADDR      =  4'h0;
parameter REG_UART_CONTROL_ADDR     =  4'h1;
parameter REG_UART_WRITE_FIFO_ADDR  =  4'h2;
parameter REG_UART_READ_FIFO_ADDR   =  4'h3;
