`include "test_base.sv"
`include "test_packet_fix.sv"
