parameter   REG_FRAC_CTRL_STATUS        = 4'h0 ;
parameter   REG_FRAC_CX_7_0_ADDR        = 4'h1 ;
parameter   REG_FRAC_CX_15_8_ADDR       = 4'h2 ;
parameter   REG_FRAC_CX_23_16_ADDR      = 4'h3 ;
parameter   REG_FRAC_CX_31_24_ADDR      = 4'h4 ;
parameter   REG_FRAC_CY_7_0_ADDR        = 4'h5 ;
parameter   REG_FRAC_CY_15_8_ADDR       = 4'h6 ;
parameter   REG_FRAC_CY_23_16_ADDR      = 4'h7 ;
parameter   REG_FRAC_CY_31_24_ADDR      = 4'h8 ;
parameter   REG_FRAC_MAX_ITER_LOW_ADDR  = 4'h9 ;
parameter   REG_FRAC_MAX_ITER_HIGH_ADDR = 4'ha ;
parameter   REG_FRAC_PY_7_0_ADDR        = 4'hb ;
parameter   REG_FRAC_PY_15_8_ADDR       = 4'hc ;
parameter   REG_FRAC_PX_7_0_ADDR        = 4'hd ;
parameter   REG_FRAC_PX_15_8_ADDR       = 4'he ;
