


// Instantiate the module
clock_gen instance_name (
    .CLKIN_IN(CLKIN_IN), 
    .CLKDV_OUT(CLKDV_OUT), 
    .CLKFX_OUT(CLKFX_OUT), 
    .CLKIN_IBUFG_OUT(CLKIN_IBUFG_OUT), 
    .CLK0_OUT(CLK0_OUT), 
    .CLK2X_OUT(CLK2X_OUT), 
    .LOCKED_OUT(LOCKED_OUT)
    );


