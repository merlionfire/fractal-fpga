module ascii_font16X8 (
   input  wire         clk,
   input  wire [10:0]  font_bitmap_addr,
   output wire  [7:0]  font_bitmap_byte 
);

// Simulation model 
/* 
   reg [7:0]   bitmap_reg [ 0 : 2047 ] ; 
   reg         font_bitmap_byte_r ; 

   assign   font_bitmap_byte =  font_bitmap_byte_r ;   
   initial begin 
      $readmemh("../rtl/ascii_font16x8.mem", bitmap_reg, 0, 2047 ) ;    
   end 

   always @( posedge clk ) begin  
      font_bitmap_byte_r <= bitmap_reg[ font_bitmap_addr] ;  
   end 
*/
   // 128 ascii chars' 16X8 font bitmap  
   RAMB16_S9 #(
    .INIT    ( 9'h000 ),     
    .INIT_00 ( 256'h00_00_00_00_7e_81_81_99_bd_81_81_a5_81_7e_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00 ),
    .INIT_01 ( 256'h00_00_00_00_10_38_7c_fe_fe_fe_fe_6c_00_00_00_00_00_00_00_00_7e_ff_ff_e7_c3_ff_ff_db_ff_7e_00_00 ),
    .INIT_02 ( 256'h00_00_00_00_3c_18_18_e7_e7_e7_3c_3c_18_00_00_00_00_00_00_00_00_10_38_7c_fe_7c_38_10_00_00_00_00 ),
    .INIT_03 ( 256'h00_00_00_00_00_00_18_3c_3c_18_00_00_00_00_00_00_00_00_00_00_3c_18_18_7e_ff_ff_7e_3c_18_00_00_00 ),
    .INIT_04 ( 256'h00_00_00_00_00_3c_66_42_42_66_3c_00_00_00_00_00_ff_ff_ff_ff_ff_ff_e7_c3_c3_e7_ff_ff_ff_ff_ff_ff ),
    .INIT_05 ( 256'h00_00_00_00_78_cc_cc_cc_cc_78_32_1a_0e_1e_00_00_ff_ff_ff_ff_ff_c3_99_bd_bd_99_c3_ff_ff_ff_ff_ff ),
    .INIT_06 ( 256'h00_00_00_00_e0_f0_70_30_30_30_30_3f_33_3f_00_00_00_00_00_00_18_18_7e_18_3c_66_66_66_66_3c_00_00 ),
    .INIT_07 ( 256'h00_00_00_00_18_18_db_3c_e7_3c_db_18_18_00_00_00_00_00_00_c0_e6_e7_67_63_63_63_63_7f_63_7f_00_00 ),
    .INIT_08 ( 256'h00_00_00_00_02_06_0e_1e_3e_fe_3e_1e_0e_06_02_00_00_00_00_00_80_c0_e0_f0_f8_fe_f8_f0_e0_c0_80_00 ),
    .INIT_09 ( 256'h00_00_00_00_66_66_00_66_66_66_66_66_66_66_00_00_00_00_00_00_00_18_3c_7e_18_18_18_7e_3c_18_00_00 ),
    .INIT_0A ( 256'h00_00_00_7c_c6_0c_38_6c_c6_c6_6c_38_60_c6_7c_00_00_00_00_00_1b_1b_1b_1b_1b_7b_db_db_db_7f_00_00 ),
    .INIT_0B ( 256'h00_00_00_00_7e_18_3c_7e_18_18_18_7e_3c_18_00_00_00_00_00_00_fe_fe_fe_fe_00_00_00_00_00_00_00_00 ),
    .INIT_0C ( 256'h00_00_00_00_18_3c_7e_18_18_18_18_18_18_18_00_00_00_00_00_00_18_18_18_18_18_18_18_7e_3c_18_00_00 ),
    .INIT_0D ( 256'h00_00_00_00_00_00_30_60_fe_60_30_00_00_00_00_00_00_00_00_00_00_00_18_0c_fe_0c_18_00_00_00_00_00 ),
    .INIT_0E ( 256'h00_00_00_00_00_00_28_6c_fe_6c_28_00_00_00_00_00_00_00_00_00_00_00_fe_c0_c0_c0_00_00_00_00_00_00 ),
    .INIT_0F ( 256'h00_00_00_00_00_10_38_38_7c_7c_fe_fe_00_00_00_00_00_00_00_00_00_fe_fe_7c_7c_38_38_10_00_00_00_00 ),
    .INIT_10 ( 256'h00_00_00_00_18_18_00_18_18_18_3c_3c_3c_18_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00 ),
    .INIT_11 ( 256'h00_00_00_00_6c_6c_fe_6c_6c_6c_fe_6c_6c_00_00_00_00_00_00_00_00_00_00_00_00_00_00_24_66_66_66_00 ),
    .INIT_12 ( 256'h00_00_00_00_86_c6_60_30_18_0c_c6_c2_00_00_00_00_00_00_18_18_7c_c6_86_06_06_7c_c0_c2_c6_7c_18_18 ),
    .INIT_13 ( 256'h00_00_00_00_00_00_00_00_00_00_00_60_30_30_30_00_00_00_00_00_76_cc_cc_cc_dc_76_38_6c_6c_38_00_00 ),
    .INIT_14 ( 256'h00_00_00_00_30_18_0c_0c_0c_0c_0c_0c_18_30_00_00_00_00_00_00_0c_18_30_30_30_30_30_30_18_0c_00_00 ),
    .INIT_15 ( 256'h00_00_00_00_00_00_18_18_7e_18_18_00_00_00_00_00_00_00_00_00_00_00_66_3c_ff_3c_66_00_00_00_00_00 ),
    .INIT_16 ( 256'h00_00_00_00_00_00_00_00_fe_00_00_00_00_00_00_00_00_00_00_30_18_18_18_00_00_00_00_00_00_00_00_00 ),
    .INIT_17 ( 256'h00_00_00_00_80_c0_60_30_18_0c_06_02_00_00_00_00_00_00_00_00_18_18_00_00_00_00_00_00_00_00_00_00 ),
    .INIT_18 ( 256'h00_00_00_00_7e_18_18_18_18_18_18_78_38_18_00_00_00_00_00_00_38_6c_c6_c6_d6_d6_c6_c6_6c_38_00_00 ),
    .INIT_19 ( 256'h00_00_00_00_7c_c6_06_06_06_3c_06_06_c6_7c_00_00_00_00_00_00_fe_c6_c0_60_30_18_0c_06_c6_7c_00_00 ),
    .INIT_1A ( 256'h00_00_00_00_7c_c6_06_06_06_fc_c0_c0_c0_fe_00_00_00_00_00_00_1e_0c_0c_0c_fe_cc_6c_3c_1c_0c_00_00 ),
    .INIT_1B ( 256'h00_00_00_00_30_30_30_30_18_0c_06_06_c6_fe_00_00_00_00_00_00_7c_c6_c6_c6_c6_fc_c0_c0_60_38_00_00 ),
    .INIT_1C ( 256'h00_00_00_00_78_0c_06_06_06_7e_c6_c6_c6_7c_00_00_00_00_00_00_7c_c6_c6_c6_c6_7c_c6_c6_c6_7c_00_00 ),
    .INIT_1D ( 256'h00_00_00_00_30_18_18_00_00_00_18_18_00_00_00_00_00_00_00_00_00_18_18_00_00_00_18_18_00_00_00_00 ),
    .INIT_1E ( 256'h00_00_00_00_00_00_00_7e_00_00_7e_00_00_00_00_00_00_00_00_00_06_0c_18_30_60_30_18_0c_06_00_00_00 ),
    .INIT_1F ( 256'h00_00_00_00_18_18_00_18_18_18_0c_c6_c6_7c_00_00_00_00_00_00_60_30_18_0c_06_0c_18_30_60_00_00_00 ),
    .INIT_20 ( 256'h00_00_00_00_c6_c6_c6_c6_fe_c6_c6_6c_38_10_00_00_00_00_00_00_7c_c0_dc_de_de_de_c6_c6_7c_00_00_00 ),
    .INIT_21 ( 256'h00_00_00_00_3c_66_c2_c0_c0_c0_c0_c2_66_3c_00_00_00_00_00_00_fc_66_66_66_66_7c_66_66_66_fc_00_00 ),
    .INIT_22 ( 256'h00_00_00_00_fe_66_62_60_68_78_68_62_66_fe_00_00_00_00_00_00_f8_6c_66_66_66_66_66_66_6c_f8_00_00 ),
    .INIT_23 ( 256'h00_00_00_00_3a_66_c6_c6_de_c0_c0_c2_66_3c_00_00_00_00_00_00_f0_60_60_60_68_78_68_62_66_fe_00_00 ),
    .INIT_24 ( 256'h00_00_00_00_3c_18_18_18_18_18_18_18_18_3c_00_00_00_00_00_00_c6_c6_c6_c6_c6_fe_c6_c6_c6_c6_00_00 ),
    .INIT_25 ( 256'h00_00_00_00_e6_66_66_6c_78_78_6c_66_66_e6_00_00_00_00_00_00_78_cc_cc_cc_0c_0c_0c_0c_0c_1e_00_00 ),
    .INIT_26 ( 256'h00_00_00_00_c6_c6_c6_c6_c6_d6_fe_fe_ee_c6_00_00_00_00_00_00_fe_66_62_60_60_60_60_60_60_f0_00_00 ),
    .INIT_27 ( 256'h00_00_00_00_7c_c6_c6_c6_c6_c6_c6_c6_c6_7c_00_00_00_00_00_00_c6_c6_c6_c6_ce_de_fe_f6_e6_c6_00_00 ),
    .INIT_28 ( 256'h00_00_0e_0c_7c_de_d6_c6_c6_c6_c6_c6_c6_7c_00_00_00_00_00_00_f0_60_60_60_60_7c_66_66_66_fc_00_00 ),
    .INIT_29 ( 256'h00_00_00_00_7c_c6_c6_06_0c_38_60_c6_c6_7c_00_00_00_00_00_00_e6_66_66_66_6c_7c_66_66_66_fc_00_00 ),
    .INIT_2A ( 256'h00_00_00_00_7c_c6_c6_c6_c6_c6_c6_c6_c6_c6_00_00_00_00_00_00_3c_18_18_18_18_18_18_5a_7e_7e_00_00 ),
    .INIT_2B ( 256'h00_00_00_00_6c_ee_fe_d6_d6_d6_c6_c6_c6_c6_00_00_00_00_00_00_10_38_6c_c6_c6_c6_c6_c6_c6_c6_00_00 ),
    .INIT_2C ( 256'h00_00_00_00_3c_18_18_18_18_3c_66_66_66_66_00_00_00_00_00_00_c6_c6_6c_7c_38_38_7c_6c_c6_c6_00_00 ),
    .INIT_2D ( 256'h00_00_00_00_3c_30_30_30_30_30_30_30_30_3c_00_00_00_00_00_00_fe_c6_c2_60_30_18_0c_86_c6_fe_00_00 ),
    .INIT_2E ( 256'h00_00_00_00_3c_0c_0c_0c_0c_0c_0c_0c_0c_3c_00_00_00_00_00_00_02_06_0e_1c_38_70_e0_c0_80_00_00_00 ),
    .INIT_2F ( 256'h00_00_ff_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_c6_6c_38_10 ),
    .INIT_30 ( 256'h00_00_00_00_76_cc_cc_cc_7c_0c_78_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_18_30_30 ),
    .INIT_31 ( 256'h00_00_00_00_7c_c6_c0_c0_c0_c6_7c_00_00_00_00_00_00_00_00_00_7c_66_66_66_66_6c_78_60_60_e0_00_00 ),
    .INIT_32 ( 256'h00_00_00_00_7c_c6_c0_c0_fe_c6_7c_00_00_00_00_00_00_00_00_00_76_cc_cc_cc_cc_6c_3c_0c_0c_1c_00_00 ),
    .INIT_33 ( 256'h00_78_cc_0c_7c_cc_cc_cc_cc_cc_76_00_00_00_00_00_00_00_00_00_f0_60_60_60_60_f0_60_64_6c_38_00_00 ),
    .INIT_34 ( 256'h00_00_00_00_3c_18_18_18_18_18_38_00_18_18_00_00_00_00_00_00_e6_66_66_66_66_76_6c_60_60_e0_00_00 ),
    .INIT_35 ( 256'h00_00_00_00_e6_66_6c_78_78_6c_66_60_60_e0_00_00_00_3c_66_66_06_06_06_06_06_06_0e_00_06_06_00_00 ),
    .INIT_36 ( 256'h00_00_00_00_c6_d6_d6_d6_d6_fe_ec_00_00_00_00_00_00_00_00_00_3c_18_18_18_18_18_18_18_18_38_00_00 ),
    .INIT_37 ( 256'h00_00_00_00_7c_c6_c6_c6_c6_c6_7c_00_00_00_00_00_00_00_00_00_66_66_66_66_66_66_dc_00_00_00_00_00 ),
    .INIT_38 ( 256'h00_1e_0c_0c_7c_cc_cc_cc_cc_cc_76_00_00_00_00_00_00_f0_60_60_7c_66_66_66_66_66_dc_00_00_00_00_00 ),
    .INIT_39 ( 256'h00_00_00_00_7c_c6_0c_38_60_c6_7c_00_00_00_00_00_00_00_00_00_f0_60_60_60_66_76_dc_00_00_00_00_00 ),
    .INIT_3A ( 256'h00_00_00_00_76_cc_cc_cc_cc_cc_cc_00_00_00_00_00_00_00_00_00_1c_36_30_30_30_30_fc_30_30_10_00_00 ),
    .INIT_3B ( 256'h00_00_00_00_6c_fe_d6_d6_d6_c6_c6_00_00_00_00_00_00_00_00_00_18_3c_66_66_66_66_66_00_00_00_00_00 ),
    .INIT_3C ( 256'h00_f8_0c_06_7e_c6_c6_c6_c6_c6_c6_00_00_00_00_00_00_00_00_00_c6_6c_38_38_38_6c_c6_00_00_00_00_00 ),
    .INIT_3D ( 256'h00_00_00_00_0e_18_18_18_18_70_18_18_18_0e_00_00_00_00_00_00_fe_c6_60_30_18_cc_fe_00_00_00_00_00 ),
    .INIT_3E ( 256'h00_00_00_00_70_18_18_18_18_0e_18_18_18_70_00_00_00_00_00_00_18_18_18_18_18_00_18_18_18_18_00_00 ),
    .INIT_3F ( 256'h00_00_00_00_00_fe_c6_c6_c6_6c_38_10_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_dc_76_00_00 ),
    // unused parity
    .INITP_00( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INITP_01( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INITP_02( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INITP_03( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INITP_04( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INITP_05( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INITP_06( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INITP_07( 256'h0000000000000000000000000000000000000000000000000000000000000000 )
   ) font16X8_inst (
    .DO     ( font_bitmap_byte ),
    .DOP    (                  ),
    .ADDR   ( font_bitmap_addr ),
    .CLK    ( clk              ),
    .DI     ( 8'h00            ),
    .DIP    ( 1'b0             ),
    .EN     ( 1'b1             ),
    .WE     ( 1'b0             ),
    .SSR    ( 1'b0             )
 );


endmodule   

